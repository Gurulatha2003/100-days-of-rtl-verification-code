 interface dff_if;
  logic clk;
  logic rst;
  logic din;
  logic dout;  
endinterface
